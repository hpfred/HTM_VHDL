library verilog;
use verilog.vl_types.all;
entity HTM_Core_vlg_vec_tst is
end HTM_Core_vlg_vec_tst;
