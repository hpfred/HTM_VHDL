LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY Memes IS
	PORT
	(
		tipos: IN ;
	);
END ENTITY Memes;

ARCHITECTURE  Carinhas OF Memes IS
BEGIN

END Carinhas;